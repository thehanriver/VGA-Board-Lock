module vga_display(
  input rst,
  input clk,
  input [19:0] ssd,

  output reg [2:0]R,
  output reg [2:0]G,
  output reg [1:0]B,
  output HS,
  output VS,
  output reg light
);
  
   
  wire [10:0] x, y;
  wire blank;
  wire cccc;
  
  clk_divider12 caseclock(clk, rst, cccc);
  
  vga_controller_640_60 vc(
    .rst(rst),
	 .pixel_clk(cccc),
	 .HS(HS),
	 .VS(VS),
	 .hcounter(x),
	 .vcounter(y),
	 .blank(blank)
  );
  
  wire clk_25Mhz;
  
clock_dividerVGA (
clk,rst, clk_25Mhz
);


 always @(posedge clk_25Mhz) begin
    light <= ~blank;
	end

  
  
  wire sq_C0,sq_C1,sq_C2,sq_C3,sq_L1, sq_S0, sq_S1, sq_S2, sq_S3, sq_D0, sq_D1, sq_D2, sq_D3, sq_A0, sq_A1, sq_A2, sq_A3, sq_B0, sq_B1, sq_B2, sq_B3, sq_E0, sq_E1, sq_E2, sq_E3;
  wire sq_F0, sq_F1, sq_F2, sq_F3, sq_00, sq_01, sq_02, sq_03, sq_10, sq_11, sq_12, sq_13, sq_20, sq_21, sq_22, sq_23, sq_30, sq_31, sq_32, sq_33, sq_40, sq_41, sq_42, sq_43, sq_44;
  wire sq_50, sq_51, sq_52, sq_53, sq_60, sq_61, sq_62, sq_63, sq_70, sq_71, sq_72, sq_73, sq_80, sq_81, sq_82, sq_83, sq_90, sq_91, sq_92, sq_93;
  wire sq_n3, sq_P2, sq_dash0, sq_dash1, sq_dash2;
  



assign sq_00 = (((x > 100) & (y >  75) & (x < 220) & (y < 115))||((x > 100) & (y >  410) & (x < 220) & (y < 450))||((x > 180) & (y >  75) & (x < 220) & (y < 450))||((x > 100) & (y >  75) & (x < 140) & (y < 450)))   ;  
    assign sq_01 = (((x > 260) & (y >  75) & (x < 380) & (y < 115))||((x > 260) & (y >  410) & (x < 380) & (y < 450))||((x > 340) & (y >  75) & (x < 380) & (y < 450))||((x > 260) & (y >  75) & (x < 300) & (y < 450)))   ;  
	 assign sq_02 = (((x > 420) & (y >  75) & (x < 540) & (y < 115))||((x > 420) & (y >  410) & (x < 540) & (y < 450))||((x > 500) & (y >  75) & (x < 540) & (y < 450))||((x > 420) & (y >  75) & (x < 460) & (y < 450)))   ;  
	 assign sq_03 = (((x > 580) & (y >  75) & (x < 700) & (y < 115))||((x > 580) & (y >  410) & (x < 700) & (y < 450))||((x > 660) & (y >  75) & (x < 700) & (y < 450))||((x > 580) & (y >  75) & (x < 620) & (y < 450)))   ;  
	

    assign sq_C0 = (((x > 100) & (y >  75) & (x < 220) & (y < 115))||((x > 100) & (y >  410) & (x < 220) & (y < 450))||((x > 100) & (y >  75) & (x < 140) & (y < 450)))  ;
	 assign sq_C1 = (((x > 260) & (y >  75) & (x < 380) & (y < 115))||((x > 260) & (y >  410) & (x < 380) & (y < 450))||((x > 260) & (y >  75) & (x < 300) & (y < 450)))  ;
	 assign sq_C2 = (((x > 420) & (y >  75) & (x < 540) & (y < 115))||((x > 420) & (y >  410) & (x < 540) & (y < 450))||((x > 420) & (y >  75) & (x < 460) & (y < 450)))  ;
	 assign sq_C3 = (((x > 580) & (y >  75) & (x < 700) & (y < 115))||((x > 580) & (y >  410) & (x < 700) & (y < 450))||((x > 580) & (y >  75) & (x < 620) & (y < 450)))  ;
    
	 assign sq_L1 = (((x > 260) & (y >  75) & (x < 300) & (y < 450)))||((x > 260) & (y >  75) & (x < 380) & (y < 115))  ;
    
	 
	 assign sq_S0 = (((x > 100) & (y >  75) & (x < 220) & (y < 115))||((x > 100) & (y >  410) & (x < 220) & (y < 450))||((x > 180) & (y >  75) & (x < 220) & (y < 275))||((x > 100) & (y >  275) & (x < 140) & (y < 450))||((x > 100) & (y >  235) & (x < 220) & (y < 275)))  ;
    assign sq_S1 = (((x > 260) & (y >  75) & (x < 380) & (y < 115))||((x > 260) & (y >  410) & (x < 380) & (y < 450))||((x > 340) & (y >  75) & (x < 380) & (y < 275))||((x > 260) & (y >  275) & (x < 300) & (y < 450))||((x > 260) & (y >  235) & (x < 380) & (y < 275)))  ;
	 assign sq_S2 = (((x > 420) & (y >  75) & (x < 540) & (y < 115))||((x > 420) & (y >  410) & (x < 540) & (y < 450))||((x > 500) & (y >  75) & (x < 540) & (y < 275))||((x > 420) & (y >  275) & (x < 460) & (y < 450))||((x > 420) & (y >  235) & (x < 540) & (y < 275)))  ;
	 assign sq_S3 = (((x > 580) & (y >  75) & (x < 700) & (y < 115))||((x > 580) & (y >  410) & (x < 700) & (y < 450))||((x > 660) & (y >  75) & (x < 700) & (y < 275))||((x > 580) & (y >  275) & (x < 620) & (y < 450))||((x > 560) & (y >  235) & (x < 700) & (y < 275)))  ;
	 
	 
	 
	 assign sq_D0 = (((x > 100) & (y >  75) & (x < 220) & (y < 115))||((x > 180) & (y >  75) & (x < 220) & (y < 450))||((x > 100) & (y >  235) & (x < 220) & (y < 275))||((x > 100) & (y >  75) & (x < 140) & (y < 235)))   ;
	 assign sq_D1 = (((x > 260) & (y >  75) & (x < 380) & (y < 115))||((x > 340) & (y >  75) & (x < 380) & (y < 450))||((x > 260) & (y >  235) & (x < 380) & (y < 275))||((x > 260) & (y >  75) & (x < 300) & (y < 235)))   ;
	 assign sq_D2 = (((x > 420) & (y >  75) & (x < 540) & (y < 115))||((x > 500) & (y >  75) & (x < 540) & (y < 450))||((x > 420) & (y >  235) & (x < 540) & (y < 275))||((x > 420) & (y >  75) & (x < 460) & (y < 235)))   ;
	 assign sq_D3 = (((x > 580) & (y >  75) & (x < 700) & (y < 115))||((x > 660) & (y >  75) & (x < 700) & (y < 450))||((x > 580) & (y >  235) & (x < 700) & (y < 275))||((x > 580) & (y >  75) & (x < 620) & (y < 235)))   ;
	 
	 
	 
	 
	 assign sq_90 = (((x > 100) & (y >  410) & (x < 220) & (y < 450))||((x > 180) & (y >  75) & (x < 220) & (y < 450))||((x > 100) & (y >  235) & (x < 220) & (y < 275))||((x > 100) & (y >  235) & (x < 140) & (y < 450)))   ;  
	 assign sq_91 = (((x > 260) & (y >  410) & (x < 380) & (y < 450))||((x > 340) & (y >  75) & (x < 380) & (y < 450))||((x > 260) & (y >  235) & (x < 380) & (y < 275))||((x > 260) & (y >  235) & (x < 300) & (y < 450)))   ;
	 assign sq_92 = (((x > 420) & (y >  410) & (x < 540) & (y < 450))||((x > 500) & (y >  75) & (x < 540) & (y < 450))||((x > 440) & (y >  235) & (x < 540) & (y < 275))||((x > 420) & (y >  235) & (x < 460) & (y < 450)))   ;
	 assign sq_93 = (((x > 580) & (y >  410) & (x < 700) & (y < 450))||((x > 660) & (y >  75) & (x < 700) & (y < 450))||((x > 620) & (y >  235) & (x < 700) & (y < 275))||((x > 580) & (y >  235) & (x < 620) & (y < 450)))   ;
	 
	 
	 
	 assign sq_80 = (((x > 100) & (y >  75) & (x < 220) & (y < 115))||((x > 100) & (y >  410) & (x < 220) & (y < 450))||((x > 180) & (y >  75) & (x < 220) & (y < 450))||((x > 100) & (y >  235) & (x < 220) & (y < 275))||((x > 100) & (y >  75) & (x < 140) & (y < 450)))   ;
	 assign sq_81 = (((x > 260) & (y >  75) & (x < 380) & (y < 115))||((x > 260) & (y >  410) & (x < 380) & (y < 450))||((x > 340) & (y >  75) & (x < 380) & (y < 450))||((x > 260) & (y >  235) & (x < 380) & (y < 275))||((x > 260) & (y >  75) & (x < 300) & (y < 450)))   ;
	 assign sq_82 = (((x > 420) & (y >  75) & (x < 540) & (y < 115))||((x > 420) & (y >  410) & (x < 540) & (y < 450))||((x > 500) & (y >  75) & (x < 540) & (y < 450))||((x > 420) & (y >  235) & (x < 540) & (y < 275))||((x > 420) & (y >  75) & (x < 460) & (y < 450)))   ;
	 assign sq_83 = (((x > 580) & (y >  75) & (x < 700) & (y < 115))||((x > 580) & (y >  410) & (x < 700) & (y < 450))||((x > 660) & (y >  75) & (x < 700) & (y < 450))||((x > 580) & (y >  235) & (x < 700) & (y < 275))||((x > 580) & (y >  75) & (x < 620) & (y < 450)))   ;
	 
	 
	 
    assign sq_70 = (((x > 100) & (y >  410) & (x < 220) & (y < 450))||((x > 180) & (y >  75) & (x < 220) & (y < 450))) ;
	 assign sq_71 = (((x > 260) & (y >  410) & (x < 380) & (y < 450))||((x > 340) & (y >  75) & (x < 380) & (y < 450))) ;
	 assign sq_72 = (((x > 420) & (y >  410) & (x < 540) & (y < 450))||((x > 500) & (y >  75) & (x < 540) & (y < 450))) ;
	 assign sq_73 = (((x > 580) & (y >  410) & (x < 700) & (y < 450))||((x > 660) & (y >  75) & (x < 700) & (y < 450))) ;
	 
	 
	 
	 assign sq_60 = (((x > 100) & (y  >  75) & (x < 220) & (y < 115))||((x > 100) & (y >  410) & (x < 220) & (y < 450))||((x > 180) & (y >  75) & (x < 220) & (y < 275))||((x > 100) & (y >  275) & (x < 140) & (y < 450))||((x > 100) & (y >  235) & (x < 220) & (y < 275)))  ;
	 assign sq_61 = (((x > 260) & (y  >  75) & (x < 380) & (y < 115))||((x > 260) & (y >  410) & (x < 380) & (y < 450))||((x > 340) & (y >  75) & (x < 380) & (y < 275))||((x > 260) & (y >  275) & (x < 300) & (y < 450))||((x > 260) & (y >  235) & (x < 380) & (y < 275)))  ;
	 assign sq_62 = (((x > 420) & (y  >  75) & (x < 540) & (y < 115))||((x > 420) & (y >  410) & (x < 540) & (y < 450))||((x > 500) & (y >  75) & (x < 540) & (y < 275))||((x > 420) & (y >  275) & (x < 460) & (y < 450))||((x > 420) & (y >  235) & (x < 540) & (y < 275)))  ;
	 assign sq_63 = (((x > 580) & (y  >  75) & (x < 700) & (y < 115))||((x > 580) & (y >  410) & (x < 700) & (y < 450))||((x > 660) & (y >  75) & (x < 700) & (y < 275))||((x > 580) & (y >  275) & (x < 620) & (y < 450))||((x > 580) & (y >  235) & (x < 700) & (y < 275)))  ;
	 
	 
	 
	 assign sq_50 = (((x > 100) & (y >  75) & (x < 220) & (y < 115))||((x > 100) & (y >  410) & (x < 220) & (y < 450))||((x > 180) & (y >  75) & (x < 220) & (y < 275))||((x > 100) & (y >  275) & (x < 140) & (y < 450))||((x > 100) & (y >  235) & (x < 220) & (y < 275)))  ;
    assign sq_51 = (((x > 260) & (y >  75) & (x < 380) & (y < 115))||((x > 260) & (y >  410) & (x < 380) & (y < 450))||((x > 340) & (y >  75) & (x < 380) & (y < 275))||((x > 260) & (y >  275) & (x < 300) & (y < 450))||((x > 260) & (y >  235) & (x < 380) & (y < 275)))  ;
	 assign sq_52 = (((x > 420) & (y >  75) & (x < 540) & (y < 115))||((x > 420) & (y >  410) & (x < 540) & (y < 450))||((x > 500) & (y >  75) & (x < 540) & (y < 275))||((x > 420) & (y >  275) & (x < 460) & (y < 450))||((x > 420) & (y >  235) & (x < 540) & (y < 275)))  ;
	 assign sq_53 = (((x > 580) & (y >  75) & (x < 700) & (y < 115))||((x > 580) & (y >  410) & (x < 700) & (y < 450))||((x > 660) & (y >  75) & (x < 700) & (y < 275))||((x > 580) & (y >  275) & (x < 620) & (y < 450))||((x > 560) & (y >  235) & (x < 700) & (y < 275)))  ;
	 
	 
	 
	 assign sq_40 = (((x > 180) & (y >  75) & (x < 220) & (y < 450))||((x > 100) & (y >  275) & (x < 140) & (y < 450))||((x > 100) & (y >  235) & (x < 220) & (y < 275)))  ;
    assign sq_41 = (((x > 340) & (y >  75) & (x < 380) & (y < 450))||((x > 260) & (y >  275) & (x < 300) & (y < 450))||((x > 260) & (y >  235) & (x < 380) & (y < 275)))  ;
    assign sq_42 = (((x > 500) & (y >  75) & (x < 540) & (y < 450))||((x > 420) & (y >  275) & (x < 460) & (y < 450))||((x > 420) & (y >  235) & (x < 540) & (y < 275)))  ;
    assign sq_43 = (((x > 660) & (y >  75) & (x < 700) & (y < 450))||((x > 580) & (y >  275) & (x < 620) & (y < 450))||((x > 580) & (y >  235) & (x < 700) & (y < 275)))  ;
    
	 
	 
	 assign sq_30 = (((x > 100) & (y >  75) & (x < 220) & (y < 115))||((x > 100) & (y >  410) & (x < 220) & (y < 450))||((x > 180) & (y >  75) & (x < 220) & (y < 450))||((x > 100) & (y >  235) & (x < 220) & (y < 275)))  ; 
    assign sq_31 = (((x > 260) & (y >  75) & (x < 380) & (y < 115))||((x > 260) & (y >  410) & (x < 380) & (y < 450))||((x > 340) & (y >  75) & (x < 380) & (y < 450))||((x > 260) & (y >  235) & (x < 380) & (y < 275)))  ; 
    assign sq_32 = (((x > 420) & (y >  75) & (x < 540) & (y < 115))||((x > 420) & (y >  410) & (x < 540) & (y < 450))||((x > 500) & (y >  75) & (x < 540) & (y < 450))||((x > 420) & (y >  235) & (x < 540) & (y < 275)))  ; 
    assign sq_33 = (((x > 580) & (y >  75) & (x < 700) & (y < 115))||((x > 580) & (y >  410) & (x < 700) & (y < 450))||((x > 660) & (y >  75) & (x < 700) & (y < 450))||((x > 580) & (y >  235) & (x < 700) & (y < 275)))  ; 
    
	 
	 
	 assign sq_20 = (((x > 100) & (y >  75) & (x < 220) & (y < 115))||((x > 100) & (y >  410) & (x < 220) & (y < 450))||((x > 100) & (y >  75) & (x < 140) & (y < 275))||((x > 180) & (y >  275) & (x < 220) & (y < 450))||((x > 100) & (y >  235) & (x < 220) & (y < 275)))  ;
    assign sq_21 = (((x > 260) & (y >  75) & (x < 380) & (y < 115))||((x > 260) & (y >  410) & (x < 380) & (y < 450))||((x > 260) & (y >  75) & (x < 300) & (y < 275))||((x > 340) & (y >  275) & (x < 380) & (y < 450))||((x > 260) & (y >  235) & (x < 380) & (y < 275)))  ;
    assign sq_22 = (((x > 420) & (y >  75) & (x < 540) & (y < 115))||((x > 420) & (y >  410) & (x < 540) & (y < 450))||((x > 420) & (y >  75) & (x < 460) & (y < 275))||((x > 500) & (y >  275) & (x < 540) & (y < 450))||((x > 420) & (y >  235) & (x < 540) & (y < 275)))  ;
    assign sq_23 = (((x > 580) & (y >  75) & (x < 700) & (y < 115))||((x > 580) & (y >  410) & (x < 700) & (y < 450))||((x > 580) & (y >  75) & (x < 620) & (y < 275))||((x > 660) & (y >  275) & (x < 700) & (y < 450))||((x > 580) & (y >  235) & (x < 700) & (y < 275)))  ;
    
	 
	 
	 assign sq_10 = ((x > 180) & (y >  75) & (x < 220) & (y < 450))  ; 
	 assign sq_11 = ((x > 340) & (y >  75) & (x < 380) & (y < 450))  ; 
	 assign sq_12 = ((x > 500) & (y >  75) & (x < 540) & (y < 450))  ; 
	 assign sq_13 = ((x > 660) & (y >  75) & (x < 700) & (y < 450))  ; 
	 
 
	 
	 
	 assign sq_A0 = (((x > 100) & (y >  410) & (x < 220) & (y < 450))||((x > 180) & (y >  75) & (x < 220) & (y < 450))||((x > 100) & (y >  235) & (x < 220) & (y < 275))||((x > 100) & (y >  75) & (x < 140) & (y < 450)))  ; 
    assign sq_A1 = (((x > 260) & (y >  410) & (x < 380) & (y < 450))||((x > 340) & (y >  75) & (x < 380) & (y < 450))||((x > 260) & (y >  235) & (x < 380) & (y < 275))||((x > 260) & (y >  75) & (x < 300) & (y < 450)))  ; 
    assign sq_A2 = (((x > 420) & (y >  410) & (x < 540) & (y < 450))||((x > 500) & (y >  75) & (x < 540) & (y < 450))||((x > 420) & (y >  235) & (x < 540) & (y < 275))||((x > 420) & (y >  75) & (x < 460) & (y < 450)))  ; 
    assign sq_A3 = (((x > 580) & (y >  410) & (x < 700) & (y < 450))||((x > 660) & (y >  75) & (x < 700) & (y < 450))||((x > 580) & (y >  235) & (x < 700) & (y < 275))||((x > 580) & (y >  75) & (x < 620) & (y < 450)))  ; 
    
	 
	 
	 assign sq_B0 = (((x > 100) & (y >  75) & (x < 220) & (y < 115))||((x > 100) & (y >  75) & (x < 140) & (y < 450))||((x > 100) & (y >  235) & (x < 220) & (y < 275))||((x > 180) & (y >  75) & (x < 220) & (y < 235)))  ;
    assign sq_B1 = (((x > 260) & (y >  75) & (x < 380) & (y < 115))||((x > 260) & (y >  75) & (x < 300) & (y < 450))||((x > 260) & (y >  235) & (x < 380) & (y < 275))||((x > 340) & (y >  75) & (x < 380) & (y < 235)))  ;
    assign sq_B2 = (((x > 420) & (y >  75) & (x < 540) & (y < 115))||((x > 420) & (y >  75) & (x < 460) & (y < 450))||((x > 420) & (y >  235) & (x < 540) & (y < 275))||((x > 500) & (y >  75) & (x < 540) & (y < 235)))  ;
    assign sq_B3 = (((x > 580) & (y >  75) & (x < 700) & (y < 115))||((x > 580) & (y >  75) & (x < 620) & (y < 450))||((x > 580) & (y >  235) & (x < 700) & (y < 275))||((x > 660) & (y >  75) & (x < 700) & (y < 235))) ;
    
	 
	 assign sq_E0 = (((x > 100) & (y >  75) & (x < 220) & (y < 115))||((x > 100) & (y >  410) & (x < 220) & (y < 450))||((x > 100) & (y >  235) & (x < 220) & (y < 275))||((x > 100) & (y >  75) & (x < 140) & (y < 450)))  ;
	 assign sq_E1 = (((x > 260) & (y >  75) & (x < 380) & (y < 115))||((x > 260) & (y >  410) & (x < 380) & (y < 450))||((x > 260) & (y >  235) & (x < 380) & (y < 275))||((x > 260) & (y >  75) & (x < 300) & (y < 450))) ;
	 assign sq_E2 = (((x > 420) & (y >  75) & (x < 540) & (y < 115))||((x > 420) & (y >  410) & (x < 540) & (y < 450))||((x > 420) & (y >  235) & (x < 540) & (y < 275))||((x > 420) & (y >  75) & (x < 460) & (y < 450))) ;
	 assign sq_E3 = (((x > 580) & (y >  75) & (x < 700) & (y < 115))||((x > 580) & (y >  410) & (x < 700) & (y < 450))||((x > 580) & (y >  235) & (x < 700) & (y < 275))||((x > 580) & (y >  75) & (x < 620) & (y < 450)))  ;
	 
	 
	 assign sq_F0 = (((x > 100) & (y >  410) & (x < 220) & (y < 450))||((x > 100) & (y >  235) & (x < 220) & (y < 275))||((x > 100) & (y >  75) & (x < 140) & (y < 450)))  ;
    assign sq_F1 = (((x > 260) & (y >  410) & (x < 380) & (y < 450))||((x > 260) & (y >  235) & (x < 380) & (y < 275))||((x > 260) & (y >  75) & (x < 300) & (y < 450))) ;
    assign sq_F2 = (((x > 420) & (y >  410) & (x < 540) & (y < 450))||((x > 420) & (y >  235) & (x < 540) & (y < 275))||((x > 420) & (y >  75) & (x < 460) & (y < 450))) ;
    assign sq_F3 = (((x > 580) & (y >  410) & (x < 700) & (y < 450))||((x > 580) & (y >  235) & (x < 700) & (y < 275))||((x > 580) & (y >  75) & (x < 620) & (y < 450))) ;
    
	 
	 assign sq_dash0 = ((x > 100) & (y >  235) & (x < 220) & (y < 275)) ;
	 assign sq_dash1 = ((x > 100) & (y >  235) & (x < 220) & (y < 275)) ;
	 assign sq_dash2 = ((x > 100) & (y >  235) & (x < 220) & (y < 275));
	 
	 
	 assign sq_P1 = (((x > 260) & (y >  410) & (x < 380) & (y < 450))||((x > 340) & (y >  275) & (x < 380) & (y < 450))||((x > 260) & (y >  235) & (x < 380) & (y < 275))||((x > 260) & (y >  75) & (x < 300) & (y < 450)));
	 
    assign sq_n3 = (((x > 580) & (y >  235) & (x < 700) & (y < 275))||((x > 660) & (y >  75) & (x < 700) & (y < 235))||((x > 580) & (y >  75) & (x < 620) & (y < 235)));



 
	
	
always @(ssd) begin
	case (ssd[19:15])
	5'b00000: begin 
	if(sq_00 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b00001: begin
	if(sq_10 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b00010: begin 
	if(sq_20 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b00011: begin
	if(sq_30 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b00100: begin 
	if(sq_40 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b00101: begin
	if(sq_50 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b00110: begin 
	if(sq_60 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b00111: begin
	if(sq_70 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
 
  5'b01000: begin 
	if(sq_80 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b01001: begin
	if(sq_90 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b01010: begin 
	if(sq_A0 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b01011: begin
	if(sq_B0 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b01100: begin 
	if(sq_C0 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b01101: begin
	if(sq_D0 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b01110: begin 
	if(sq_E0 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b01111: begin
	if(sq_F0 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b10000: begin
	if(sq_C0 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b10010: begin 
	if(sq_S0 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b11111: begin
	if(sq_dash0 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  default: begin
  R = 3'b000;
  G = 3'b111;
  B = 2'b00;
  end
  endcase  
 

 
  case (ssd[14:10])
	
	5'b00000: begin 
	if(sq_01 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b00001: begin
	if(sq_11 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b00010: begin 
	if(sq_21 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b00011: begin
	if(sq_31 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b00100: begin 
	if(sq_41 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b00101: begin
	if(sq_51 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b00110: begin 
	if(sq_61 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b00111: begin
	if(sq_71 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  
  
  
  5'b01000: begin 
	if(sq_81 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b01001: begin
	if(sq_91 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b01010: begin 
	if(sq_A1 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b01011: begin
	if(sq_B1 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b01100: begin 
	if(sq_C1 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b01101: begin
	if(sq_D1 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b01110: begin 
	if(sq_E1 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b01111: begin
	if(sq_F1 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b10000: begin
	if(sq_C1 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b10010: begin 
	if(sq_S1 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b11111: begin
	if(sq_dash1 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  
  
  5'b10001: begin 
	if(sq_L1 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b10111: begin
	if(sq_P1 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  default: begin
  R = 3'b000;
  G = 3'b111;
  B = 2'b00;
  end
  endcase
  
  
  
  case (ssd[9:5])
	
	5'b00000: begin 
	if(sq_02 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b00001: begin
	if(sq_12 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b00010: begin 
	if(sq_22 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b00011: begin
	if(sq_32 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b00100: begin 
	if(sq_42 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b00101: begin
	if(sq_52 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b00110: begin 
	if(sq_62 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b00111: begin
	if(sq_72 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  
  
  
  5'b01000: begin 
	if(sq_82 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b01001: begin
	if(sq_92 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b01010: begin 
	if(sq_A2 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b01011: begin
	if(sq_B2 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b01100: begin 
	if(sq_C2 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b01101: begin
	if(sq_D2 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b01110: begin 
	if(sq_E2 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b01111: begin
	if(sq_F2 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b10000: begin
	if(sq_C2 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b10010: begin 
	if(sq_S2 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b11111: begin
	if(sq_dash2 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
 default: begin
  R = 3'b000;
  G = 3'b111;
  B = 2'b00;
  end
  endcase
  
  case (ssd[4:0])
	
	5'b00000: begin 
	if(sq_03 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b00001: begin
	if(sq_13 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b00010: begin 
	if(sq_23 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b00011: begin
	if(sq_33 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b00100: begin 
	if(sq_43 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b00101: begin
	if(sq_53 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b00110: begin 
	if(sq_63 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b00111: begin
	if(sq_73 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  
  
  
  5'b01000: begin 
	if(sq_83 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b01001: begin
	if(sq_93 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b01010: begin 
	if(sq_A3 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b01011: begin
	if(sq_B3 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b01100: begin 
	if(sq_C3 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b01101: begin
	if(sq_D3 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b01110: begin 
	if(sq_E3 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b01111: begin
	if(sq_F3 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b10000: begin
	if(sq_C3 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  
  5'b10010: begin 
	if(sq_S3 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
   
	5'b11000: begin
	if(sq_n3 == 1) begin
	R = 3'b000;
	G = 3'b111;
	B = 2'b00;
	end
  end
  default: begin
  R = 3'b000;
  G = 3'b111;
  B = 2'b00;
  end
  endcase
  end
endmodule
